`define BARREL_SHIFTER
`undef  SHIFTER
`define ACTING_LOW
`undef  ACTING_HIGH
`define CLK_INNER 50000000
`define FREQ_SHIFT 10
`define FREQ_FOR_ANODES 5000
